module example1;
    initial begin $display("Hello World"); $finish; end
endmodule

