.title KiCad schematic
J1 __J1
U1 __U1
U2 __U2
X1 __X1
.end
